magic
tech sky130A
timestamp 1759450942
<< nwell >>
rect 0 0 160 100
<< ndiff >>
rect 90 58 115 70
rect 90 42 98 58
rect 107 42 115 58
rect 90 30 115 42
<< pdiff >>
rect 30 58 60 70
rect 30 42 40 58
rect 50 42 60 58
rect 30 30 60 42
<< ndiffc >>
rect 98 42 107 58
<< pdiffc >>
rect 40 42 50 58
<< metal1 >>
rect 40 42 50 58
rect 98 42 107 58
<< end >>
